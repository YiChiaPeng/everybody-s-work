library verilog;
use verilog.vl_types.all;
entity ripple_4bit_UP_counter_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ripple_4bit_UP_counter_vlg_sample_tst;
