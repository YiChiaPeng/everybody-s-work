library verilog;
use verilog.vl_types.all;
entity ripple_DOWN_counter_vlg_vec_tst is
end ripple_DOWN_counter_vlg_vec_tst;
