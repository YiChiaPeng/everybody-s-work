library verilog;
use verilog.vl_types.all;
entity ripple_4bit_UP_counter_vlg_vec_tst is
end ripple_4bit_UP_counter_vlg_vec_tst;
