library verilog;
use verilog.vl_types.all;
entity ripple_DOWN_counter_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ripple_DOWN_counter_vlg_sample_tst;
