library verilog;
use verilog.vl_types.all;
entity sametime_counter_12bit_vlg_vec_tst is
end sametime_counter_12bit_vlg_vec_tst;
